module main

import gx

const (
	screen_height = 480
	screen_width = 640

	bg_color = gx.black
)