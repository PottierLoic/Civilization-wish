module main

import gx

const (
	// Dimensions
	screen_height = 640
	screen_width = 640
	cell_size = 20

	// Colors
	bg_color = gx.black
	desert_color = gx.yellow
	forest_color = gx.green
	sea_color = gx.blue
)