module main

struct Biome {
	name string

}

fn new_biome() Biome {
	return Biome{
		name: 'desert'
	}
}