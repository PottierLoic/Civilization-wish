module main

import gx

const (
	// Dimensions
	screen_width = 300
	screen_height = 300
	cell_size = 40

	// Colors
	bg_color = gx.black
)