module main

import gx

const (
	// Dimensions
	screen_height = 500
	screen_width = 500
	cell_size = 10

	// Colors
	bg_color = gx.black
	sand_color = gx.rgb(240, 240, 64)
	forest_color = gx.rgb(16, 160, 0)
	shallow_water_color = gx.rgb(25, 25, 150)
	deep_water_color = gx.rgb(0, 0, 128)
	grass_color = gx.rgb(50, 220, 20)
	rock_color = gx.rgb(128, 128, 128)
	snow_color = gx.rgb(255, 255, 255)

)