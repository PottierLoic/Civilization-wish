module main

struct Game {
	mut:
		world World
		players Player
}